`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    04/14/2023 
// Design Name: 
// Module Name:    DFF_INT_TEST_TOP 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module DFF_INT_TEST_TOP(
    input CLK_50M,
    input save_data_dff_pi,

    input DB_DFFQ0_1,
    input DB_DFFQ0_2,
    input DB_DFFQ0_3,
    input DB_DFFQ0_4,
    input DB_DFFQ0_5,
    input DB_DFFQ0_6,
    input DB_DFFQ0_7,
    input DB_DFFQ0_8,
    input DB_DFFQ0_9,
    input DB_DFFQ1_0,
    input DB_DFFQ1_1,
    input DB_DFFQ1_2,
    input DB_DFFQ1_3,
    input DB_DFFQ1_4,
    input DB_DFFQ1_5,
    input DB_DFFQ1_6,
    input DB_DFFQ1_7,
    input DB_DFFQ1_8,
    input DB_DFFQ1_9,

    input data_clk_dff_pi,
    output data_out_dff_pi,
);

endmodule
